* C:\Users\chinm\eSim-Workspace\inv_testing\inv_testing.cir

.include inv_A.sub
X1  in vdd out inv_A		
		
Vdd vdd 0 3.3
vd0 in 0 pulse(0 1.8 0s 0s 0s 5us 10us)

.tran 0.1us 40us

.control
run

plot V(in) 
plot V(out)

.endc
.end
