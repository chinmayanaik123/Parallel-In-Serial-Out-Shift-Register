* C:\Users\chinm\eSim-Workspace\dff_testing\dff_testing.cir

.include dff_A.sub
		
X1  din clk vdd qout dff_A		
		
		
Vdd vdd 0 3.3
vd0 din 0 pulse(0 1.8 0s 0s 0s 10us 20us)
vd1 clk 0 pulse(0 1.8 0s 0s 0s 5us 10us)
.tran 0.1us 40us

.control
run
plot V(clk)
plot V(din) 
plot V(qout)

.endc
.end